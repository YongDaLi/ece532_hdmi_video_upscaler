`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/02/2023 01:41:59 AM
// Design Name: 
// Module Name: tb_mario_processing
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module tb_mario_processing();
    chunk_input last_chunk;
    chunk_input current_chunk;
    
    chunk_output current_output_chunk;
    chunk_output next_output_chunk;
    
    
    processor p(
        .last_chunk(last_chunk),
        .current_chunk(current_chunk),
        .output_chunk_current(current_output_chunk),
        .output_chunk_next(next_output_chunk)
    );
    
    initial begin
        last_chunk = {{ { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 } }, { { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 } }, { { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'h8b, 8'h45, 8'h00 } }, { { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 }, { 8'h99, 8'h69, 8'h1a }, { 8'h8b, 8'h45, 8'h00 } }, { { 8'h8b, 8'h45, 8'h00 }, { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a } }, { { 8'h99, 8'h69, 8'h1a }, { 8'h00, 8'h00, 8'h00 }, { 8'h99, 8'h69, 8'h1a }, { 8'h00, 8'h00, 8'h00 } }, { { 8'h99, 8'h69, 8'h1a }, { 8'hff, 8'hff, 8'hff }, { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'h99, 8'h69, 8'h1a }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'h8b, 8'h45, 8'h00 }, { 8'hff, 8'hff, 8'hff }, { 8'h8b, 8'h45, 8'h00 } }, { { 8'h99, 8'h69, 8'h1a }, { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 }, { 8'h99, 8'h69, 8'h1a } }, { { 8'h8b, 8'h45, 8'h00 }, { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a } }, { { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a }, { 8'h00, 8'h00, 8'h00 } }, { { 8'h00, 8'h00, 8'h00 }, { 8'h99, 8'h69, 8'h1a }, { 8'h00, 8'h00, 8'h00 }, { 8'h00, 8'h00, 8'h00 } }, { { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a }, { 8'h00, 8'h00, 8'h00 }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'h99, 8'h69, 8'h1a }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 } }, { { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a }, { 8'h00, 8'h00, 8'hff }, { 8'hff, 8'h00, 8'h00 } }, { { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 } }, { { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 } }, { { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 } }, { { 8'h00, 8'h00, 8'hff }, { 8'hff, 8'h00, 8'h00 }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff } }, { { 8'hff, 8'h00, 8'h00 }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff } }, { { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 } }, { { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'h00, 8'h00 }, { 8'h00, 8'h00, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'h00, 8'h00, 8'hff } }, { { 8'hff, 8'hff, 8'h00 }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff } }, { { 8'h00, 8'h00, 8'hff }, { 8'hff, 8'hff, 8'h00 }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff } }, { { 8'h00, 8'h00, 8'hff }, { 8'hff, 8'h00, 8'h00 }, { 8'h00, 8'h00, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff } }, { { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'h00, 8'h00, 8'hff } }, { { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 } }, { { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 } }, { { 8'h8b, 8'h45, 8'h00 }, { 8'hff, 8'hff, 8'hff }, { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } } };
        current_chunk = {{ { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'h00, 8'h00 } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'h99, 8'h69, 8'h1a }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 } }, { { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'h8b, 8'h45, 8'h00 }, { 8'h99, 8'h69, 8'h1a } }, { { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'h99, 8'h69, 8'h1a }, { 8'h00, 8'h00, 8'h00 } }, { { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'h99, 8'h69, 8'h1a }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'h00, 8'h00 }, { 8'h99, 8'h69, 8'h1a }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 } }, { { 8'h99, 8'h69, 8'h1a }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'h8b, 8'h45, 8'h00 }, { 8'hff, 8'hff, 8'hff }, { 8'h8b, 8'h45, 8'h00 } }, { { 8'h99, 8'h69, 8'h1a }, { 8'h8b, 8'h45, 8'h00 }, { 8'h99, 8'h69, 8'h1a }, { 8'h8b, 8'h45, 8'h00 } }, { { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a }, { 8'h8b, 8'h45, 8'h00 }, { 8'h99, 8'h69, 8'h1a } }, { { 8'h99, 8'h69, 8'h1a }, { 8'h00, 8'h00, 8'h00 }, { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a } }, { { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a }, { 8'h00, 8'h00, 8'h00 }, { 8'h99, 8'h69, 8'h1a } }, { { 8'h99, 8'h69, 8'h1a }, { 8'hff, 8'h00, 8'h00 }, { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a } }, { { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'h8b, 8'h45, 8'h00 }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'h8b, 8'h45, 8'h00 }, { 8'h99, 8'h69, 8'h1a }, { 8'hff, 8'hff, 8'hff }, { 8'h99, 8'h69, 8'h1a } }, { { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a } }, { { 8'h99, 8'h69, 8'h1a }, { 8'h00, 8'h00, 8'h00 }, { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a } }, { { 8'h00, 8'h00, 8'h00 }, { 8'h00, 8'h00, 8'h00 }, { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a } }, { { 8'h00, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a } }, { { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 } }, { { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 } }, { { 8'h00, 8'h00, 8'hff }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'h00, 8'h00, 8'hff } }, { { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 } }, { { 8'h00, 8'h00, 8'hff }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'h00, 8'h00, 8'hff } }, { { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 } }, { { 8'h99, 8'h69, 8'h1a }, { 8'h99, 8'h69, 8'h1a }, { 8'hff, 8'hff, 8'hff }, { 8'h99, 8'h69, 8'h1a } }, { { 8'h99, 8'h69, 8'h1a }, { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'h00, 8'h00 }, { 8'hff, 8'h00, 8'h00 }, { 8'h00, 8'h00, 8'hff }, { 8'hff, 8'h00, 8'h00 } }, { { 8'hff, 8'h00, 8'h00 }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff } }, { { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'hff, 8'hff, 8'h00 }, { 8'h00, 8'h00, 8'hff } }, { { 8'h00, 8'h00, 8'hff }, { 8'hff, 8'hff, 8'h00 }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff } }, { { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff } }, { { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'h8b, 8'h45, 8'h00 } }, { { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 } }, { { 8'h8b, 8'h45, 8'h00 }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff } }, { { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff } }, { { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff } }, { { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'h00, 8'h00, 8'hff }, { 8'h00, 8'h00, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'h8b, 8'h45, 8'h00 }, { 8'h8b, 8'h45, 8'h00 }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'h8b, 8'h45, 8'h00 }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'h8b, 8'h45, 8'h00 }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } }, { { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff }, { 8'hff, 8'hff, 8'hff } } };
        
        $display("Last Input");
        #20 $display("%x", current_chunk);
        $display("Current Input");
        #20 $display("%x", last_chunk);
        
        $display("Current Output");
        #20 $display("%x", current_output_chunk);
        
        $display("Next Output");
        #20 $display("%x", next_output_chunk);
    end
endmodule
